// Code your testbench here
// or browse Examples

`include "params_pkg.sv"

`include "axi_uvm_pkg.sv"

`include "tb.sv"


/*! \mainpage My Personal Index Page
 *
 * \section intro_sec Introduction
 *
 * This is the introduction.
 *
 * \section install_sec Installation
 *
 * \subsection step1 Step 1: Opening the box
 *
 * etc...
 */

// Code your testbench here
// or browse Examples

`include "params_pkg.sv"

`include "axi_uvm_pkg.sv"

`include "tb.sv"

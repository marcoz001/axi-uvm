// Code your design here

`include "params_pkg.sv"

`include "axi_pkg.sv"

`include "axi_if.sv"


// Code your design here

`include "axi_pkg.sv"

`include "axim2wbsp.v"
`include "aximrd2wbsp.v"
`include "aximwr2wbsp.v"

`include "axi_if.sv"
`include "wb_if.sv"
`include "wbarbiter.v"

// Code your design here

`include "axi_pkg.sv"

`include "axi_if.sv"



package params_pkg;

  parameter AXI_ID_WIDTH   = 6;
  parameter AXI_ADDR_WIDTH = 32;
  parameter AXI_DATA_WIDTH = 32;


endpackage : params_pkg
